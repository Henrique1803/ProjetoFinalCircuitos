library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM2 is
port(
	  address: in std_logic_vector(3 downto 0);
	  output : out std_logic_vector(31 downto 0)
);
end ROM2;

architecture arc_ROM2 of ROM2 is
begin

--         HEX7      HEX6     HEX5     HEX4     HEX3     HEX2     HEX1     HEX0               round

output <= "0101"	& "1111" & "0100" & "1111"	& "0011" & "1111" & "0010" & "0001" when address = "0000" else

          "1001"	& "0000" & "1111" & "0110"	& "1111" & "0100" & "1111" & "0101" when address = "0001" else

			 "0111"	& "1011" & "1001" & "1000"	& "1111" & "1111" & "1111" & "0010" when address = "0010" else

			 "1111"	& "1111" & "1100" & "1010"	& "1111" & "0111" & "1001" & "1101" when address = "0011" else

			 "1110"	& "1111" & "1111" & "1111"	& "0010" & "1001" & "0100" & "0000" when address = "0100" else

			 "1110"	& "1101" & "1100" & "1011"	& "1010" & "1111" & "1111" & "1111" when address = "0101" else

			 "0101"	& "1001" & "1111" & "1110"	& "1111" & "1100" & "1111" & "1000" when address = "0110" else

			 "0001"	& "0010" & "1111" & "1111"	& "1111" & "0011" & "1010" & "1011" when address = "0111" else

			 "1111"	& "1000" & "1111" & "0100"	& "1111" & "0000" & "0110" & "0010" when address = "1000" else

			 "0000"	& "1111" & "1010" & "1001"	& "1111" & "1111" & "1100" & "0111" when address = "1001" else

			 "0001"	& "1001" & "1111" & "1110"	& "1111" & "0010" & "1111" & "1101" when address = "1010" else

			 "1000"	& "1010" & "1011" & "1101"	& "1111" & "1111" & "1001" & "1111" when address = "1011" else

			 "1111"	& "1111" & "1111" & "0111"	& "0110" & "0101" & "1001" & "0000" when address = "1100" else

			 "1010"	& "1111" & "1011" & "1100"	& "0011" & "1111" & "1111" & "1101" when address = "1101" else

			 "1001"	& "1000" & "0111" & "1111"	& "0010" & "1111" & "1111" & "0000" when address = "1110" else

			 "0001"	& "1100" & "1111" & "0111"	& "1111" & "1111" & "1011" & "0011";

end arc_ROM2;